package config is

    constant N : integer := 2;
    constant M : integer := 2;
    constant NODES : integer := 4;

end package ; -- aegean_def
