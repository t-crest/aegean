library ieee;
use ieee.std_logic_1164.all;

package ocp_config is

    constant BURST_ADDR_WIDTH : integer := 27;

end package ; -- ocp_config
