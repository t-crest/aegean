package config is

    constant N : integer := 2;
    constant M : integer := 2;

end package ; -- aegean_def
