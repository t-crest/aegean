-- -----------------------------------------------------------------------------
--  Title      :  4 phase latch controllers with reset.
--
--  Notes      :  To avoid optimization of the synthesis tool
--                (Xilinx ISE), this code forces the values of the LUT.
--                This description is specifically written for the Xilinx
--                Spartan-IIE FPGA. It should synthesize on Xilinx Virtex, Virtex-E,
--                Virtex-II, Virtex-II Pro, Virtex-II Pro X, Spartan-II,
--                Spartan-IIE, and Spartan-3, but this has not been tested.
--
--                By using the UNISIM lib, ModelSim or any other VHDL simulator
--                can be used to verify the funcionality of the design.
--
--  Developer  :  Mikkel Stensgaard  -- s001434@student.dtu.dk
--
--  Revision   :  1.0    09-06-04     Initial version
-- -----------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

LIBRARY UNISIM;
USE UNISIM.Vcomponents.all;

entity AS_bd_4p_LatchController_ud is
Generic (reset_value : bit := '0');
Port ( req_in:  in  std_logic;
      ack_in:  out std_logic;
      req_out: out std_logic;
      ack_out: in  std_logic;
      reset:   in  std_logic; --active low
      lt:      out std_logic);--active high
end entity;

architecture un_decoupled of AS_bd_4p_LatchController_ud is
-----------------------
-- XILINX COMPONENTS --
-----------------------
-- 4-Bit Look-Up-Table with Local Output
component LUT4_L
generic (INIT : bit_vector(15 downto 0));
port (
      I0 : in  std_ulogic;
      I1 : in  std_ulogic;
      I2 : in  std_ulogic;
      I3 : in  std_ulogic;
      lO : out std_ulogic);
end component;

----------------------------------------------------
--# Generated by petrify 4.0 (compiled 22-Dec-98 at 8:44 AM)
--INORDER = Rin Aout Lt Rout Ain;
--OUTORDER = [Lt] [Rout] [Ain];
--[Lt] = Rout;
--[Rout] = Rin (Rout + Aout') + Aout' Rout;
--[Ain] = Lt;
--
-- the logical equation defining the C element is:
-- Rout = reset(Rin Rout + Rin Aout' + Aout' Rout)

-- Constant using the generic "reset_value"
constant rv : bit := reset_value;
constant reset_vector : bit_vector(7 downto 0) := rv&rv&rv&rv&rv&rv&rv&rv;

-- Internal signals
signal s_out : std_logic;

begin

--------------
-- Rout = reset( Rin Rout + Rin Aout' + Aout' Rout)
--------------
latch_controller: LUT4_L
generic map (INIT => "10110010"&reset_vector)
port map (I0 => req_in, I1 => ack_out, I2 => s_out, I3 => reset, LO => s_out);

--------------
-- Connect the outputs to the correct signals
--------------
req_out <= s_out;
lt <= s_out;
ack_in <= s_out;

end architecture; --ud




